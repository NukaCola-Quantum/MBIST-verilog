`timescale 1ns / 1ps
/*
//////////////////////////////////////////////////////////////////////////////////
//   Copyright 2013 - 2019 Yang Song
//   E-mail: googotohell@gmail.com
//
//   Licensed under the Apache License, Version 2.0 (the "License");
//   you may not use this file except in compliance with the License.
//   You may obtain a copy of the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in writing, software
//   distributed under the License is distributed on an "AS IS" BASIS,
//   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//   See the License for the specific language governing permissions and
//   limitations under the License.
*/
//////////////////////////////////////////////////////////////////////////////////
// Company: <-blank->
// Engineer: Yang Song
// 
// Create Date:		10:21:31 01/03/2014 
// Design Name:		FW-MBIST
// Module Name:		MBIST_TAP_interface
// Project Name: 	<-blank->
// Target Devices:	[VirtexII-FG256]
// Tool versions:  ISE 10.1(x64) QuestaSim 10.x(x64)
// Description: 
// The module designs to meet generic DFT and jtag test. It works on scan mode
// and could bypass on other ways.
// 
// Dependencies: MBIST_CONTROLLER.v, MBIST_comparator_WF.v
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/*
module MBIST_TAP_interface (
	algsel_scan_in, algsel_scan_en, algsel_scan_out, algsel_clock
	);

	input algsel_scan_in;
	input algsel_scan_en;
	input algsel_clock;
	output algsel_scan_out;
	
endmodule
*/
