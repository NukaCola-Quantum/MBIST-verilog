`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: <-blank->
// Engineer: Yang Song
// 
// Create Date:		10:21:31 01/03/2014 
// Design Name:		MBIST_diagnostics
// Module Name:		MBIST_diagnostics
// Project Name: 	<-blank->
// Target Devices:	[VirtexII-FG256]
// Tool versions:  ISE 10.1(x64) QuestaSim 10.x(x64)
// Description: 
// (MBIST_diagnostics block should exactly locate fail bits position and output
// other details about errors. It needs to custom depend on UUT.)
// 
// Dependencies: None
//
// Revision:
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/*
module MBIST_diagnostics (
	diag_scan_in, diag_clk, rst_h, hold_l, debugz, diag_scan_out, diag_monitor
	);
	
	input diag_scan_in;
	input diag_clk;
	input rst_h;
	input hold_l;
	input debugz;
	output diag_scan_out;
	output diag_monitor;
	
	
endmodule
*/
