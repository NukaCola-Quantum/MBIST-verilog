`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: <-blank->
// Engineer: Yang Song
// 
// Create Date:		10:21:31 01/03/2014 
// Design Name:		MBIST_TAP_interface
// Module Name:		MBIST_TAP_interface
// Project Name: 	<-blank->
// Target Devices:	[VirtexII-FG256]
// Tool versions:  ISE 10.1(x64) QuestaSim 10.x(x64)
// Description: 
// The module designs to meet generic DFT and jtag test. It works on scan mode
// and could bypass on other ways.
// 
// Dependencies: MBIST_CONTROLLER.v, MBIST_comparator_WF.v
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/*
module MBIST_TAP_interface (
	algsel_scan_in, algsel_scan_en, algsel_scan_out, algsel_clock
	);

	input algsel_scan_in;
	input algsel_scan_en;
	input algsel_clock;
	output algsel_scan_out;
	
endmodule
*/
