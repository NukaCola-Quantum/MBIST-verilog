`timescale 1ns / 1ps
/*
//////////////////////////////////////////////////////////////////////////////////
//   Copyright 2013 - 2019 Yang Song
//   E-mail: googotohell@gmail.com
//
//   Licensed under the Apache License, Version 2.0 (the "License");
//   you may not use this file except in compliance with the License.
//   You may obtain a copy of the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in writing, software
//   distributed under the License is distributed on an "AS IS" BASIS,
//   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//   See the License for the specific language governing permissions and
//   limitations under the License.
*/
//////////////////////////////////////////////////////////////////////////////////
// Company: <-blank->
// Engineer: Yang Song
// 
// Create Date:		10:21:31 01/03/2014 
// Design Name:		FW-MBIST
// Module Name:		MBIST_diagnostics
// Project Name: 	<-blank->
// Target Devices:	[VirtexII-FG256]
// Tool versions:  ISE 10.1(x64) QuestaSim 10.x(x64)
// Description: 
// (MBIST_diagnostics block should exactly locate fail bits position and output
// other details about errors. It needs to custom depend on UUT.)
// 
// Dependencies: None
//
// Revision:
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
/*
module MBIST_diagnostics (
	diag_scan_in, diag_clk, rst_h, hold_l, debugz, diag_scan_out, diag_monitor
	);
	
	input diag_scan_in;
	input diag_clk;
	input rst_h;
	input hold_l;
	input debugz;
	output diag_scan_out;
	output diag_monitor;
	
	
endmodule
*/
